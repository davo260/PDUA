LIBRARY	IEEE;
USE		IEEE.STD_LOGIC_1164.ALL;
USE 		IEEE.NUMERIC_STD.ALL;

ENTITY	dq_ALU	IS
	GENERIC(	DATA_WIDTH	:	INTEGER	:=	8);
				
	PORT(
				mdr_alu_n		:	IN		 STD_LOGIC;
				
				B_Bus_IN		   :	IN		 STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
				
				dq_ALU			:	INOUT  STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
		  );

END dq_ALU;

ARCHITECTURE RTL OF	dq_ALU	IS

BEGIN
	dq_ALU	<= (B_Bus_IN) WHEN mdr_alu_n='0' ELSE "ZZZZZZZZ";

END ARCHITECTURE;